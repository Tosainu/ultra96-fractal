module fractal_axi #(
  // Width of S_AXI data bus
  parameter integer S_AXI_DATA_WIDTH = 32,
  // Width of S_AXI address bus
  parameter integer S_AXI_ADDR_WIDTH = 4,
  parameter integer REGISTER_WIDTH = (2**S_AXI_ADDR_WIDTH) * 8
) (
  output reg [REGISTER_WIDTH - 1:0] registers,

  // Global Clock Signal
  input wire  S_AXI_ACLK,
  // Global Reset Signal. This Signal is Active LOW
  input wire  S_AXI_ARESETN,
  // Write address (issued by master, acceped by Slave)
  input wire [S_AXI_ADDR_WIDTH-1 : 0] S_AXI_AWADDR,
  // Write channel Protection type. This signal indicates the
      // privilege and security level of the transaction, and whether
      // the transaction is a data access or an instruction access.
  input wire [2 : 0] S_AXI_AWPROT,
  // Write address valid. This signal indicates that the master signaling
      // valid write address and control information.
  input wire  S_AXI_AWVALID,
  // Write address ready. This signal indicates that the slave is ready
      // to accept an address and associated control signals.
  output wire  S_AXI_AWREADY,
  // Write data (issued by master, acceped by Slave)
  input wire [S_AXI_DATA_WIDTH-1 : 0] S_AXI_WDATA,
  // Write strobes. This signal indicates which byte lanes hold
      // valid data. There is one write strobe bit for each eight
      // bits of the write data bus.
  input wire [(S_AXI_DATA_WIDTH/8)-1 : 0] S_AXI_WSTRB,
  // Write valid. This signal indicates that valid write
      // data and strobes are available.
  input wire  S_AXI_WVALID,
  // Write ready. This signal indicates that the slave
      // can accept the write data.
  output wire  S_AXI_WREADY,
  // Write response. This signal indicates the status
      // of the write transaction.
  output wire [1 : 0] S_AXI_BRESP,
  // Write response valid. This signal indicates that the channel
      // is signaling a valid write response.
  output wire  S_AXI_BVALID,
  // Response ready. This signal indicates that the master
      // can accept a write response.
  input wire  S_AXI_BREADY,
  // Read address (issued by master, acceped by Slave)
  input wire [S_AXI_ADDR_WIDTH-1 : 0] S_AXI_ARADDR,
  // Protection type. This signal indicates the privilege
      // and security level of the transaction, and whether the
      // transaction is a data access or an instruction access.
  input wire [2 : 0] S_AXI_ARPROT,
  // Read address valid. This signal indicates that the channel
      // is signaling valid read address and control information.
  input wire  S_AXI_ARVALID,
  // Read address ready. This signal indicates that the slave is
      // ready to accept an address and associated control signals.
  output wire  S_AXI_ARREADY,
  // Read data (issued by slave)
  output wire [S_AXI_DATA_WIDTH-1 : 0] S_AXI_RDATA,
  // Read response. This signal indicates the status of the
      // read transfer.
  output wire [1 : 0] S_AXI_RRESP,
  // Read valid. This signal indicates that the channel is
      // signaling the required read data.
  output wire  S_AXI_RVALID,
  // Read ready. This signal indicates that the master can
      // accept the read data and response information.
  input wire  S_AXI_RREADY
);

// AXI4LITE signals
reg [S_AXI_ADDR_WIDTH-1 : 0]  axi_awaddr;
reg   axi_awready;
reg   axi_wready;
reg [1 : 0]   axi_bresp;
reg   axi_bvalid;
reg [S_AXI_ADDR_WIDTH-1 : 0]  axi_araddr;
reg   axi_arready;
reg [S_AXI_DATA_WIDTH-1 : 0]  axi_rdata;
reg [1 : 0]   axi_rresp;
reg   axi_rvalid;

wire   slv_reg_rden;
wire   slv_reg_wren;
reg [S_AXI_DATA_WIDTH-1:0]   reg_data_out;
reg  aw_en;

wire [S_AXI_DATA_WIDTH-1:0] wsrtb_mask;
genvar byte_index;
for (byte_index = 0; byte_index < (S_AXI_DATA_WIDTH / 8); byte_index = byte_index + 1) begin
  assign wsrtb_mask[(byte_index * 8)+:8] = {8{S_AXI_WSTRB[byte_index]}};
end

localparam integer ADDR_LSB = (S_AXI_DATA_WIDTH / 32) + 1;

function [S_AXI_ADDR_WIDTH - 1:0] align_reg_addr;
  input [S_AXI_ADDR_WIDTH - 1:0] addr;
  align_reg_addr = {addr[S_AXI_ADDR_WIDTH - 1:ADDR_LSB], {ADDR_LSB{1'b0}}};
endfunction

wire [S_AXI_ADDR_WIDTH - 1:0] aligned_awaddr = align_reg_addr(axi_awaddr);
wire [S_AXI_ADDR_WIDTH - 1:0] aligned_araddr = align_reg_addr(axi_araddr);

// I/O Connections assignments
assign S_AXI_AWREADY = axi_awready;
assign S_AXI_WREADY  = axi_wready;
assign S_AXI_BRESP   = axi_bresp;
assign S_AXI_BVALID  = axi_bvalid;
assign S_AXI_ARREADY = axi_arready;
assign S_AXI_RDATA   = axi_rdata;
assign S_AXI_RRESP   = axi_rresp;
assign S_AXI_RVALID  = axi_rvalid;

// Implement axi_awready generation
// axi_awready is asserted for one S_AXI_ACLK clock cycle when both
// S_AXI_AWVALID and S_AXI_WVALID are asserted. axi_awready is
// de-asserted when reset is low.
always @(posedge S_AXI_ACLK) begin
  if (S_AXI_ARESETN == 1'b0) begin
    axi_awready <= 1'b0;
    aw_en <= 1'b1;
  end
  else begin
    if (~axi_awready && S_AXI_AWVALID && S_AXI_WVALID && aw_en) begin
      // slave is ready to accept write address when
      // there is a valid write address and write data
      // on the write address and data bus. This design
      // expects no outstanding transactions.
      axi_awready <= 1'b1;
      aw_en <= 1'b0;
    end
    else if (S_AXI_BREADY && axi_bvalid) begin
      aw_en <= 1'b1;
      axi_awready <= 1'b0;
    end
    else begin
        axi_awready <= 1'b0;
    end
  end
end

// Implement axi_awaddr latching
// This process is used to latch the address when both
// S_AXI_AWVALID and S_AXI_WVALID are valid.
always @(posedge S_AXI_ACLK) begin
  if (S_AXI_ARESETN == 1'b0)
    begin
      axi_awaddr <= 0;
    end
  else
    begin
      if (~axi_awready && S_AXI_AWVALID && S_AXI_WVALID && aw_en)
        begin
          // Write Address latching
          axi_awaddr <= S_AXI_AWADDR;
        end
    end
end

// Implement axi_wready generation
// axi_wready is asserted for one S_AXI_ACLK clock cycle when both
// S_AXI_AWVALID and S_AXI_WVALID are asserted. axi_wready is
// de-asserted when reset is low.
always @(posedge S_AXI_ACLK) begin
  if (S_AXI_ARESETN == 1'b0) begin
    axi_wready <= 1'b0;
  end
  else begin
    if (~axi_wready && S_AXI_WVALID && S_AXI_AWVALID && aw_en ) begin
      // slave is ready to accept write data when
      // there is a valid write address and write data
      // on the write address and data bus. This design
      // expects no outstanding transactions.
      axi_wready <= 1'b1;
    end
    else begin
      axi_wready <= 1'b0;
    end
  end
end

// Implement memory mapped register select and write logic generation
// The write data is accepted and written to memory mapped registers when
// axi_awready, S_AXI_WVALID, axi_wready and S_AXI_WVALID are asserted. Write strobes are used to
// select byte enables of slave registers while writing.
// These registers are cleared when reset (active low) is applied.
// Slave register write enable is asserted when valid address and data are available
// and the slave is ready to accept the write address and write data.
assign slv_reg_wren = axi_wready && S_AXI_WVALID && axi_awready && S_AXI_AWVALID;

always @(posedge S_AXI_ACLK) begin
  if (S_AXI_ARESETN == 1'b0)
    registers <= 'h0;
  else
    if (slv_reg_wren)
      registers[{aligned_awaddr, 3'b000}+:S_AXI_DATA_WIDTH] <= (S_AXI_WDATA & wsrtb_mask) | (registers[{aligned_awaddr, 3'b000}+:S_AXI_DATA_WIDTH] & ~wsrtb_mask);
end

// Implement write response logic generation
// The write response and response valid signals are asserted by the slave
// when axi_wready, S_AXI_WVALID, axi_wready and S_AXI_WVALID are asserted.
// This marks the acceptance of address and indicates the status of
// write transaction.

always @(posedge S_AXI_ACLK) begin
  if (S_AXI_ARESETN == 1'b0) begin
    axi_bvalid  <= 0;
    axi_bresp   <= 2'b0;
  end
  else begin
    if (axi_awready && S_AXI_AWVALID && ~axi_bvalid && axi_wready && S_AXI_WVALID) begin
      // indicates a valid write response is available
      axi_bvalid <= 1'b1;
      axi_bresp  <= 2'b0; // 'OKAY' response
    end                   // work error responses in future
    else begin
      if (S_AXI_BREADY && axi_bvalid) begin
        //check if bready is asserted while bvalid is high)
        //(there is a possibility that bready is always asserted high)
        axi_bvalid <= 1'b0;
      end
    end
  end
end

// Implement axi_arready generation
// axi_arready is asserted for one S_AXI_ACLK clock cycle when
// S_AXI_ARVALID is asserted. axi_awready is
// de-asserted when reset (active low) is asserted.
// The read address is also latched when S_AXI_ARVALID is
// asserted. axi_araddr is reset to zero on reset assertion.
always @(posedge S_AXI_ACLK) begin
  if (S_AXI_ARESETN == 1'b0) begin
    axi_arready <= 1'b0;
    axi_araddr  <= 32'b0;
  end
  else begin
    if (~axi_arready && S_AXI_ARVALID) begin
      // indicates that the slave has acceped the valid read address
      axi_arready <= 1'b1;
      // Read address latching
      axi_araddr  <= S_AXI_ARADDR;
    end
    else begin
      axi_arready <= 1'b0;
    end
  end
end

// Implement axi_arvalid generation
// axi_rvalid is asserted for one S_AXI_ACLK clock cycle when both
// S_AXI_ARVALID and axi_arready are asserted. The slave registers
// data are available on the axi_rdata bus at this instance. The
// assertion of axi_rvalid marks the validity of read data on the
// bus and axi_rresp indicates the status of read transaction.axi_rvalid
// is deasserted on reset (active low). axi_rresp and axi_rdata are
// cleared to zero on reset (active low).
always @(posedge S_AXI_ACLK) begin
  if (S_AXI_ARESETN == 1'b0) begin
    axi_rvalid <= 0;
    axi_rresp  <= 0;
  end
  else begin
    if (axi_arready && S_AXI_ARVALID && ~axi_rvalid) begin
      // Valid read data is available at the read data bus
      axi_rvalid <= 1'b1;
      axi_rresp  <= 2'b0; // 'OKAY' response
    end
    else if (axi_rvalid && S_AXI_RREADY) begin
      // Read data is accepted by the master
      axi_rvalid <= 1'b0;
    end
  end
end

// Implement memory mapped register select and read logic generation
// Slave register read enable is asserted when valid address is available
// and the slave is ready to accept the read address.
assign slv_reg_rden = axi_arready & S_AXI_ARVALID & ~axi_rvalid;
always @(*) begin
  reg_data_out <= registers[{aligned_araddr, 3'b000}+:S_AXI_DATA_WIDTH];
end

// Output register or memory read data
always @(posedge S_AXI_ACLK) begin
  if (S_AXI_ARESETN == 1'b0) begin
    axi_rdata  <= 0;
  end
  else begin
    // When there is a valid read address (S_AXI_ARVALID) with
    // acceptance of read address by the slave (axi_arready),
    // output the read dada
    if (slv_reg_rden) begin
      axi_rdata <= reg_data_out;     // register read data
    end
  end
end

endmodule
